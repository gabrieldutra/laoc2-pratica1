library verilog;
use verilog.vl_types.all;
entity pratica1 is
    port(
        clock           : in     vl_logic
    );
end pratica1;
